library verilog;
use verilog.vl_types.all;
entity one_pulse is
    port(
        clk             : in     vl_logic;
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end one_pulse;
