library verilog;
use verilog.vl_types.all;
entity note_player_tb_v is
    generic(
        delay           : integer := 10
    );
end note_player_tb_v;
