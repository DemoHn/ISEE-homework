library verilog;
use verilog.vl_types.all;
entity sine_reader_tb_v is
    generic(
        delay           : integer := 10
    );
end sine_reader_tb_v;
