library verilog;
use verilog.vl_types.all;
entity mcu_tb_v is
    generic(
        delay           : integer := 10
    );
end mcu_tb_v;
