module sine_rom (
  clk, dout, addr,i
);
	input clk;
	input i;
	output [15 : 0] dout;
	input [9 : 0] addr;

	wire [15:0] memory [1023:0];
	reg [15:0] dout;

	always @(posedge clk)
		begin
			if(i)
				dout = ~memory[addr];
			else
				dout = memory[addr];
		end
   

assign memory[	0	]=	16'd	0            ;
assign memory[	1	]=	16'd	50           ;
assign memory[	2	]=	16'd	101     	;
assign memory[	3	]=	16'd	151     	;
assign memory[	4	]=	16'd	201     	;
assign memory[	5	]=	16'd	251     	;
assign memory[	6	]=	16'd	302     	;
assign memory[	7	]=	16'd	352     	;
assign memory[	8	]=	16'd	402     	;
assign memory[	9	]=	16'd	452     	;
assign memory[	10	]=	16'd	503     	;
assign memory[	11	]=	16'd	553     	;
assign memory[	12	]=	16'd	603          ;
assign memory[	13	]=	16'd	653     	;
assign memory[	14	]=	16'd	704          ;
assign memory[	15	]=	16'd	754     	;
assign memory[	16	]=	16'd	804     	;
assign memory[	17	]=	16'd	854     	;
assign memory[	18	]=	16'd	905     	;
assign memory[	19	]=	16'd	955     	;
assign memory[	20	]=	16'd	1005    	;
assign memory[	21	]=	16'd	1055    	;
assign memory[	22	]=	16'd	1106    	;
assign memory[	23	]=	16'd	1156    	;
assign memory[	24	]=	16'd	1206    	;
assign memory[	25	]=	16'd	1256         ;
assign memory[	26	]=	16'd	1307    	;
assign memory[	27	]=	16'd	1357    	;
assign memory[	28	]=	16'd	1407    	;
assign memory[	29	]=	16'd	1457    	;
assign memory[	30	]=	16'd	1507    	;
assign memory[	31	]=	16'd	1558    	;
assign memory[	32	]=	16'd	1608    	;
assign memory[	33	]=	16'd	1658    	;
assign memory[	34	]=	16'd	1708    	;
assign memory[	35	]=	16'd	1758    	;
assign memory[	36	]=	16'd	1809    	;
assign memory[	37	]=	16'd	1859    	;
assign memory[	38	]=	16'd	1909    	;
assign memory[	39	]=	16'd	1959    	;
assign memory[	40	]=	16'd	2009    	;
assign memory[	41	]=	16'd	2059    	;
assign memory[	42	]=	16'd	2110    	;
assign memory[	43	]=	16'd	2160    	;
assign memory[	44	]=	16'd	2210         ;
assign memory[	45	]=	16'd	2260    	;
assign memory[	46	]=	16'd	2310    	;
assign memory[	47	]=	16'd	2360    	;
assign memory[	48	]=	16'd	2410    	;
assign memory[	49	]=	16'd	2461    	;
assign memory[	50	]=	16'd	2511    	;
assign memory[	51	]=	16'd	2561    	;
assign memory[	52	]=	16'd	2611    	;
assign memory[	53	]=	16'd	2661    	;
assign memory[	54	]=	16'd	2711    	;
assign memory[	55	]=	16'd	2761    	;
assign memory[	56	]=	16'd	2811    	;
assign memory[	57	]=	16'd	2861    	;
assign memory[	58	]=	16'd	2911    	;
assign memory[	59	]=	16'd	2962    	;
assign memory[	60	]=	16'd	3012    	;
assign memory[	61	]=	16'd	3062    	;
assign memory[	62	]=	16'd	3112    	;
assign memory[	63	]=	16'd	3162    	;
assign memory[	64	]=	16'd	3212         ;
assign memory[	65	]=	16'd	3262    	;
assign memory[	66	]=	16'd	3312    	;
assign memory[	67	]=	16'd	3362    	;
assign memory[	68	]=	16'd	3412    	;
assign memory[	69	]=	16'd	3462    	;
assign memory[	70	]=	16'd	3512    	;
assign memory[	71	]=	16'd	3562    	;
assign memory[	72	]=	16'd	3612    	;
assign memory[	73	]=	16'd	3662    	;
assign memory[	74	]=	16'd	3712    	;
assign memory[	75	]=	16'd	3761    	;
assign memory[	76	]=	16'd	3811    	;
assign memory[	77	]=	16'd	3861    	;
assign memory[	78	]=	16'd	3911    	;
assign memory[	79	]=	16'd	3961    	;
assign memory[	80	]=	16'd	4011    	;
assign memory[	81	]=	16'd	4061    	;
assign memory[	82	]=	16'd	4111    	;
assign memory[	83	]=	16'd	4161    	;
assign memory[	84	]=	16'd	4210    	;
assign memory[	85	]=	16'd	4260    	;
assign memory[	86	]=	16'd	4310    	;
assign memory[	87	]=	16'd	4360    	;
assign memory[	88	]=	16'd	4410    	;
assign memory[	89	]=	16'd	4460    	;
assign memory[	90	]=	16'd	4509    	;
assign memory[	91	]=	16'd	4559    	;
assign memory[	92	]=	16'd	4609    	;
assign memory[	93	]=	16'd	4659    	;
assign memory[	94	]=	16'd	4708    	;
assign memory[	95	]=	16'd	4758    	;
assign memory[	96	]=	16'd	4808    	;
assign memory[	97	]=	16'd	4858    	;
assign memory[	98	]=	16'd	4907    	;
assign memory[	99	]=	16'd	4957    	;
assign memory[	100	]=	16'd	5007 		;
assign memory[	101	]=	16'd	5056 		;
assign memory[	102	]=	16'd	5106 		;
assign memory[	103	]=	16'd	5156 		;
assign memory[	104	]=	16'd	5205 		;
assign memory[	105	]=	16'd	5255 		;
assign memory[	106	]=	16'd	5305 		;
assign memory[	107	]=	16'd	5354 		;
assign memory[	108	]=	16'd	5404 	     ;
assign memory[	109	]=	16'd	5453 		;
assign memory[	110	]=	16'd	5503 		;
assign memory[	111	]=	16'd	5552 		;
assign memory[	112	]=	16'd	5602 		;
assign memory[	113	]=	16'd	5651 		;
assign memory[	114	]=	16'd	5701 		;
assign memory[	115	]=	16'd	5750 		;
assign memory[	116	]=	16'd	5800 	     ;
assign memory[	117	]=	16'd	5849 		;
assign memory[	118	]=	16'd	5899 		;
assign memory[	119	]=	16'd	5948 		;
assign memory[	120	]=	16'd	5998 		;
assign memory[	121	]=	16'd	6047 		;
assign memory[	122	]=	16'd	6096 		;
assign memory[	123	]=	16'd	6146 		;
assign memory[	124	]=	16'd	6195 		;
assign memory[	125	]=	16'd	6245 		;
assign memory[	126	]=	16'd	6294 		;
assign memory[	127	]=	16'd	6343 		;
assign memory[	128	]=	16'd	6393 		;
assign memory[	129	]=	16'd	6442 		;
assign memory[	130	]=	16'd	6491 		;
assign memory[	131	]=	16'd	6540 		;
assign memory[	132	]=	16'd	6590 		;
assign memory[	133	]=	16'd	6639 		;
assign memory[	134	]=	16'd	6688 		;
assign memory[	135	]=	16'd	6737 		;
assign memory[	136	]=	16'd	6786 		;
assign memory[	137	]=	16'd	6836 		;
assign memory[	138	]=	16'd	6885 		;
assign memory[	139	]=	16'd	6934 		;
assign memory[	140	]=	16'd	6983 	     ;
assign memory[	141	]=	16'd	7032 		;
assign memory[	142	]=	16'd	7081 		;
assign memory[	143	]=	16'd	7130 		;
assign memory[	144	]=	16'd	7179 	     ;
assign memory[	145	]=	16'd	7228 	     ;
assign memory[	146	]=	16'd	7277 		;
assign memory[	147	]=	16'd	7326 		;
assign memory[	148	]=	16'd	7375 		;
assign memory[	149	]=	16'd	7424 		;
assign memory[	150	]=	16'd	7473 		;
assign memory[	151	]=	16'd	7522 		;
assign memory[	152	]=	16'd	7571 		;
assign memory[	153	]=	16'd	7620 		;
assign memory[	154	]=	16'd	7669 		;
assign memory[	155	]=	16'd	7718 		;
assign memory[	156	]=	16'd	7767 		;
assign memory[	157	]=	16'd	7815 		;
assign memory[	158	]=	16'd	7864 		;
assign memory[	159	]=	16'd	7913 		;
assign memory[	160	]=	16'd	7962 	     ;
assign memory[	161	]=	16'd	8010 		;
assign memory[	162	]=	16'd	8059 	     ;
assign memory[	163	]=	16'd	8108 		;
assign memory[	164	]=	16'd	8157 		;
assign memory[	165	]=	16'd	8205 		;
assign memory[	166	]=	16'd	8254 		;
assign memory[	167	]=	16'd	8303 		;
assign memory[	168	]=	16'd	8351 	     ;
assign memory[	169	]=	16'd	8400 		;
assign memory[	170	]=	16'd	8448 		;
assign memory[	171	]=	16'd	8497 		;
assign memory[	172	]=	16'd	8545 		;
assign memory[	173	]=	16'd	8594 		;
assign memory[	174	]=	16'd	8642 		;
assign memory[	175	]=	16'd	8691 	     ;
assign memory[	176	]=	16'd	8739 		;
assign memory[	177	]=	16'd	8788 		;
assign memory[	178	]=	16'd	8836 		;
assign memory[	179	]=	16'd	8885 	     ;
assign memory[	180	]=	16'd	8933 		;
assign memory[	181	]=	16'd	8981 	     ;
assign memory[	182	]=	16'd	9030 		;
assign memory[	183	]=	16'd	9078 	     ;
assign memory[	184	]=	16'd	9126 		;
assign memory[	185	]=	16'd	9175 		;
assign memory[	186	]=	16'd	9223 		;
assign memory[	187	]=	16'd	9271 	     ;
assign memory[	188	]=	16'd	9319 		;
assign memory[	189	]=	16'd	9367 		;
assign memory[	190	]=	16'd	9416 	     ;
assign memory[	191	]=	16'd	9464 		;
assign memory[	192	]=	16'd	9512 		;
assign memory[	193	]=	16'd	9560 		;
assign memory[	194	]=	16'd	9608 		;
assign memory[	195	]=	16'd	9656 		;
assign memory[	196	]=	16'd	9704 		;
assign memory[	197	]=	16'd	9752 		;
assign memory[	198	]=	16'd	9800 		;
assign memory[	199	]=	16'd	9848 		;
assign memory[	200	]=	16'd	9896 		;
assign memory[	201	]=	16'd	9944 		;
assign memory[	202	]=	16'd	9992 	     ;
assign memory[	203	]=	16'd	10039		;
assign memory[	204	]=	16'd	10087	     ;
assign memory[	205	]=	16'd	10135	     ;
assign memory[	206	]=	16'd	10183		;
assign memory[	207	]=	16'd	10231		;
assign memory[	208	]=	16'd	10278	     ;
assign memory[	209	]=	16'd	10326		;
assign memory[	210	]=	16'd	10374		;
assign memory[	211	]=	16'd	10421		;
assign memory[	212	]=	16'd	10469		;
assign memory[	213	]=	16'd	10517		;
assign memory[	214	]=	16'd	10564		;
assign memory[	215	]=	16'd	10612		;
assign memory[	216	]=	16'd	10659		;
assign memory[	217	]=	16'd	10707		;
assign memory[	218	]=	16'd	10754		;
assign memory[	219	]=	16'd	10802		;
assign memory[	220	]=	16'd	10849		;
assign memory[	221	]=	16'd	10897	     ;
assign memory[	222	]=	16'd	10944		;
assign memory[	223	]=	16'd	10992		;
assign memory[	224	]=	16'd	11039		;
assign memory[	225	]=	16'd	11086		;
assign memory[	226	]=	16'd	11133		;
assign memory[	227	]=	16'd	11181		;
assign memory[	228	]=	16'd	11228		;
assign memory[	229	]=	16'd	11275		;
assign memory[	230	]=	16'd	11322		;
assign memory[	231	]=	16'd	11370		;
assign memory[	232	]=	16'd	11417	     ;
assign memory[	233	]=	16'd	11464	     ;
assign memory[	234	]=	16'd	11511		;
assign memory[	235	]=	16'd	11558		;
assign memory[	236	]=	16'd	11605		;
assign memory[	237	]=	16'd	11652		;
assign memory[	238	]=	16'd	11699		;
assign memory[	239	]=	16'd	11746		;
assign memory[	240	]=	16'd	11793		;
assign memory[	241	]=	16'd	11840		;
assign memory[	242	]=	16'd	11886		;
assign memory[	243	]=	16'd	11933	     ;
assign memory[	244	]=	16'd	11980		;
assign memory[	245	]=	16'd	12027		;
assign memory[	246	]=	16'd	12074	     ;
assign memory[	247	]=	16'd	12120		;
assign memory[	248	]=	16'd	12167		;
assign memory[	249	]=	16'd	12214		;
assign memory[	250	]=	16'd	12260		;
assign memory[	251	]=	16'd	12307		;
assign memory[	252	]=	16'd	12353	     ;
assign memory[	253	]=	16'd	12400		;
assign memory[	254	]=	16'd	12446		;
assign memory[	255	]=	16'd	12493		;
assign memory[	256	]=	16'd	12539		;
assign memory[	257	]=	16'd	12586		;
assign memory[	258	]=	16'd	12632		;
assign memory[	259	]=	16'd	12679		;
assign memory[	260	]=	16'd	12725		;
assign memory[	261	]=	16'd	12771		;
assign memory[	262	]=	16'd	12817		;
assign memory[	263	]=	16'd	12864		;
assign memory[	264	]=	16'd	12910	     ;
assign memory[	265	]=	16'd	12956		;
assign memory[	266	]=	16'd	13002		;
assign memory[	267	]=	16'd	13048		;
assign memory[	268	]=	16'd	13094	     ;
assign memory[	269	]=	16'd	13141		;
assign memory[	270	]=	16'd	13187		;
assign memory[	271	]=	16'd	13233		;
assign memory[	272	]=	16'd	13279		;
assign memory[	273	]=	16'd	13324		;
assign memory[	274	]=	16'd	13370		;
assign memory[	275	]=	16'd	13416		;
assign memory[	276	]=	16'd	13462		;
assign memory[	277	]=	16'd	13508		;
assign memory[	278	]=	16'd	13554		;
assign memory[	279	]=	16'd	13599		;
assign memory[	280	]=	16'd	13645	     ;
assign memory[	281	]=	16'd	13691		;
assign memory[	282	]=	16'd	13736		;
assign memory[	283	]=	16'd	13782		;
assign memory[	284	]=	16'd	13828		;
assign memory[	285	]=	16'd	13873		;
assign memory[	286	]=	16'd	13919		;
assign memory[	287	]=	16'd	13964		;
assign memory[	288	]=	16'd	14010		;
assign memory[	289	]=	16'd	14055		;
assign memory[	290	]=	16'd	14101		;
assign memory[	291	]=	16'd	14146		;
assign memory[	292	]=	16'd	14191		;
assign memory[	293	]=	16'd	14236		;
assign memory[	294	]=	16'd	14282	     ;
assign memory[	295	]=	16'd	14327		;
assign memory[	296	]=	16'd	14372		;
assign memory[	297	]=	16'd	14417		;
assign memory[	298	]=	16'd	14462		;
assign memory[	299	]=	16'd	14507		;
assign memory[	300	]=	16'd	14553		;
assign memory[	301	]=	16'd	14598		;
assign memory[	302	]=	16'd	14643	     ;
assign memory[	303	]=	16'd	14688		;
assign memory[	304	]=	16'd	14732	     ;
assign memory[	305	]=	16'd	14777		;
assign memory[	306	]=	16'd	14822		;
assign memory[	307	]=	16'd	14867		;
assign memory[	308	]=	16'd	14912		;
assign memory[	309	]=	16'd	14956		;
assign memory[	310	]=	16'd	15001		;
assign memory[	311	]=	16'd	15046		;
assign memory[	312	]=	16'd	15090		;
assign memory[	313	]=	16'd	15135		;
assign memory[	314	]=	16'd	15180		;
assign memory[	315	]=	16'd	15224		;
assign memory[	316	]=	16'd	15269		;
assign memory[	317	]=	16'd	15313		;
assign memory[	318	]=	16'd	15358		;
assign memory[	319	]=	16'd	15402		;
assign memory[	320	]=	16'd	15446		;
assign memory[	321	]=	16'd	15491		;
assign memory[	322	]=	16'd	15535		;
assign memory[	323	]=	16'd	15579		;
assign memory[	324	]=	16'd	15623	     ;
assign memory[	325	]=	16'd	15667		;
assign memory[	326	]=	16'd	15712		;
assign memory[	327	]=	16'd	15756		;
assign memory[	328	]=	16'd	15800		;
assign memory[	329	]=	16'd	15844		;
assign memory[	330	]=	16'd	15888		;
assign memory[	331	]=	16'd	15932		;
assign memory[	332	]=	16'd	15976	     ;
assign memory[	333	]=	16'd	16019		;
assign memory[	334	]=	16'd	16063		;
assign memory[	335	]=	16'd	16107		;
assign memory[	336	]=	16'd	16151		;
assign memory[	337	]=	16'd	16195		;
assign memory[	338	]=	16'd	16238		;
assign memory[	339	]=	16'd	16282		;
assign memory[	340	]=	16'd	16325		;
assign memory[	341	]=	16'd	16369		;
assign memory[	342	]=	16'd	16413		;
assign memory[	343	]=	16'd	16456		;
assign memory[	344	]=	16'd	16499		;
assign memory[	345	]=	16'd	16543		;
assign memory[	346	]=	16'd	16586		;
assign memory[	347	]=	16'd	16630		;
assign memory[	348	]=	16'd	16673		;
assign memory[	349	]=	16'd	16716		;
assign memory[	350	]=	16'd	16759	     ;
assign memory[	351	]=	16'd	16802		;
assign memory[	352	]=	16'd	16846		;
assign memory[	353	]=	16'd	16889		;
assign memory[	354	]=	16'd	16932		;
assign memory[	355	]=	16'd	16975		;
assign memory[	356	]=	16'd	17018	     ;
assign memory[	357	]=	16'd	17061		;
assign memory[	358	]=	16'd	17104		;
assign memory[	359	]=	16'd	17146		;
assign memory[	360	]=	16'd	17189		;
assign memory[	361	]=	16'd	17232		;
assign memory[	362	]=	16'd	17275		;
assign memory[	363	]=	16'd	17317		;
assign memory[	364	]=	16'd	17360		;
assign memory[	365	]=	16'd	17403		;
assign memory[	366	]=	16'd	17445		;
assign memory[	367	]=	16'd	17488		;
assign memory[	368	]=	16'd	17530	     ;
assign memory[	369	]=	16'd	17573		;
assign memory[	370	]=	16'd	17615		;
assign memory[	371	]=	16'd	17657		;
assign memory[	372	]=	16'd	17700		;
assign memory[	373	]=	16'd	17742		;
assign memory[	374	]=	16'd	17784		;
assign memory[	375	]=	16'd	17827		;
assign memory[	376	]=	16'd	17869		;
assign memory[	377	]=	16'd	17911		;
assign memory[	378	]=	16'd	17953		;
assign memory[	379	]=	16'd	17995		;
assign memory[	380	]=	16'd	18037		;
assign memory[	381	]=	16'd	18079		;
assign memory[	382	]=	16'd	18121		;
assign memory[	383	]=	16'd	18163		;
assign memory[	384	]=	16'd	18204		;
assign memory[	385	]=	16'd	18246		;
assign memory[	386	]=	16'd	18288		;
assign memory[	387	]=	16'd	18330		;
assign memory[	388	]=	16'd	18371		;
assign memory[	389	]=	16'd	18413		;
assign memory[	390	]=	16'd	18454		;
assign memory[	391	]=	16'd	18496		;
assign memory[	392	]=	16'd	18537		;
assign memory[	393	]=	16'd	18579		;
assign memory[	394	]=	16'd	18620		;
assign memory[	395	]=	16'd	18661		;
assign memory[	396	]=	16'd	18703		;
assign memory[	397	]=	16'd	18744		;
assign memory[	398	]=	16'd	18785		;
assign memory[	399	]=	16'd	18826		;
assign memory[	400	]=	16'd	18868		;
assign memory[	401	]=	16'd	18909		;
assign memory[	402	]=	16'd	18950		;
assign memory[	403	]=	16'd	18991		;
assign memory[	404	]=	16'd	19032		;
assign memory[	405	]=	16'd	19072	     ;
assign memory[	406	]=	16'd	19113		;
assign memory[	407	]=	16'd	19154		;
assign memory[	408	]=	16'd	19195		;
assign memory[	409	]=	16'd	19236		;
assign memory[	410	]=	16'd	19276		;
assign memory[	411	]=	16'd	19317		;
assign memory[	412	]=	16'd	19357		;
assign memory[	413	]=	16'd	19398		;
assign memory[	414	]=	16'd	19438		;
assign memory[	415	]=	16'd	19479		;
assign memory[	416	]=	16'd	19519		;
assign memory[	417	]=	16'd	19560		;
assign memory[	418	]=	16'd	19600		;
assign memory[	419	]=	16'd	19640		;
assign memory[	420	]=	16'd	19680		;
assign memory[	421	]=	16'd	19721		;
assign memory[	422	]=	16'd	19761		;
assign memory[	423	]=	16'd	19801		;
assign memory[	424	]=	16'd	19841		;
assign memory[	425	]=	16'd	19881		;
assign memory[	426	]=	16'd	19921		;
assign memory[	427	]=	16'd	19961		;
assign memory[	428	]=	16'd	20000		;
assign memory[	429	]=	16'd	20040		;
assign memory[	430	]=	16'd	20080		;
assign memory[	431	]=	16'd	20120		;
assign memory[	432	]=	16'd	20159		;
assign memory[	433	]=	16'd	20199		;
assign memory[	434	]=	16'd	20238		;
assign memory[	435	]=	16'd	20278		;
assign memory[	436	]=	16'd	20317		;
assign memory[	437	]=	16'd	20357		;
assign memory[	438	]=	16'd	20396		;
assign memory[	439	]=	16'd	20436		;
assign memory[	440	]=	16'd	20475		;
assign memory[	441	]=	16'd	20514		;
assign memory[	442	]=	16'd	20553		;
assign memory[	443	]=	16'd	20592		;
assign memory[	444	]=	16'd	20631		;
assign memory[	445	]=	16'd	20670	     ;
assign memory[	446	]=	16'd	20709		;
assign memory[	447	]=	16'd	20748		;
assign memory[	448	]=	16'd	20787		;
assign memory[	449	]=	16'd	20826	     ;
assign memory[	450	]=	16'd	20865		;
assign memory[	451	]=	16'd	20904		;
assign memory[	452	]=	16'd	20942		;
assign memory[	453	]=	16'd	20981		;
assign memory[	454	]=	16'd	21019		;
assign memory[	455	]=	16'd	21058		;
assign memory[	456	]=	16'd	21096		;
assign memory[	457	]=	16'd	21135		;
assign memory[	458	]=	16'd	21173		;
assign memory[	459	]=	16'd	21212		;
assign memory[	460	]=	16'd	21250		;
assign memory[	461	]=	16'd	21288		;
assign memory[	462	]=	16'd	21326		;
assign memory[	463	]=	16'd	21364		;
assign memory[	464	]=	16'd	21403		;
assign memory[	465	]=	16'd	21441		;
assign memory[	466	]=	16'd	21479		;
assign memory[	467	]=	16'd	21516		;
assign memory[	468	]=	16'd	21554		;
assign memory[	469	]=	16'd	21592		;
assign memory[	470	]=	16'd	21630		;
assign memory[	471	]=	16'd	21668		;
assign memory[	472	]=	16'd	21705		;
assign memory[	473	]=	16'd	21743		;
assign memory[	474	]=	16'd	21781		;
assign memory[	475	]=	16'd	21818		;
assign memory[	476	]=	16'd	21856		;
assign memory[	477	]=	16'd	21893		;
assign memory[	478	]=	16'd	21930		;
assign memory[	479	]=	16'd	21968	     ;
assign memory[	480	]=	16'd	22005		;
assign memory[	481	]=	16'd	22042		;
assign memory[	482	]=	16'd	22079	     ;
assign memory[	483	]=	16'd	22116		;
assign memory[	484	]=	16'd	22154		;
assign memory[	485	]=	16'd	22191	     ;
assign memory[	486	]=	16'd	22227		;
assign memory[	487	]=	16'd	22264	     ;
assign memory[	488	]=	16'd	22301		;
assign memory[	489	]=	16'd	22338		;
assign memory[	490	]=	16'd	22375		;
assign memory[	491	]=	16'd	22411		;
assign memory[	492	]=	16'd	22448		;
assign memory[	493	]=	16'd	22485		;
assign memory[	494	]=	16'd	22521		;
assign memory[	495	]=	16'd	22558		;
assign memory[	496	]=	16'd	22594		;
assign memory[	497	]=	16'd	22631		;
assign memory[	498	]=	16'd	22667		;
assign memory[	499	]=	16'd	22703		;
assign memory[	500	]=	16'd	22739		;
assign memory[	501	]=	16'd	22776		;
assign memory[	502	]=	16'd	22812		;
assign memory[	503	]=	16'd	22848		;
assign memory[	504	]=	16'd	22884		;
assign memory[	505	]=	16'd	22920		;
assign memory[	506	]=	16'd	22956		;
assign memory[	507	]=	16'd	22991		;
assign memory[	508	]=	16'd	23027		;
assign memory[	509	]=	16'd	23063		;
assign memory[	510	]=	16'd	23099	     ;
assign memory[	511	]=	16'd	23134		;
assign memory[	512	]=	16'd	23170		;
assign memory[	513	]=	16'd	23205		;
assign memory[	514	]=	16'd	23241		;
assign memory[	515	]=	16'd	23276		;
assign memory[	516	]=	16'd	23311		;
assign memory[	517	]=	16'd	23347		;
assign memory[	518	]=	16'd	23382		;
assign memory[	519	]=	16'd	23417		;
assign memory[	520	]=	16'd	23452		;
assign memory[	521	]=	16'd	23487		;
assign memory[	522	]=	16'd	23522		;
assign memory[	523	]=	16'd	23557		;
assign memory[	524	]=	16'd	23592		;
assign memory[	525	]=	16'd	23627		;
assign memory[	526	]=	16'd	23662		;
assign memory[	527	]=	16'd	23697		;
assign memory[	528	]=	16'd	23731		;
assign memory[	529	]=	16'd	23766		;
assign memory[	530	]=	16'd	23801		;
assign memory[	531	]=	16'd	23835		;
assign memory[	532	]=	16'd	23870	     ;
assign memory[	533	]=	16'd	23904		;
assign memory[	534	]=	16'd	23938		;
assign memory[	535	]=	16'd	23973		;
assign memory[	536	]=	16'd	24007		;
assign memory[	537	]=	16'd	24041		;
assign memory[	538	]=	16'd	24075		;
assign memory[	539	]=	16'd	24109		;
assign memory[	540	]=	16'd	24143		;
assign memory[	541	]=	16'd	24177		;
assign memory[	542	]=	16'd	24211		;
assign memory[	543	]=	16'd	24245		;
assign memory[	544	]=	16'd	24279		;
assign memory[	545	]=	16'd	24312		;
assign memory[	546	]=	16'd	24346		;
assign memory[	547	]=	16'd	24380		;
assign memory[	548	]=	16'd	24413		;
assign memory[	549	]=	16'd	24447		;
assign memory[	550	]=	16'd	24480		;
assign memory[	551	]=	16'd	24514	     ;
assign memory[	552	]=	16'd	24547		;
assign memory[	553	]=	16'd	24580		;
assign memory[	554	]=	16'd	24613		;
assign memory[	555	]=	16'd	24647	     ;
assign memory[	556	]=	16'd	24680		;
assign memory[	557	]=	16'd	24713		;
assign memory[	558	]=	16'd	24746		;
assign memory[	559	]=	16'd	24779		;
assign memory[	560	]=	16'd	24811		;
assign memory[	561	]=	16'd	24844	     ;
assign memory[	562	]=	16'd	24877		;
assign memory[	563	]=	16'd	24910		;
assign memory[	564	]=	16'd	24942		;
assign memory[	565	]=	16'd	24975		;
assign memory[	566	]=	16'd	25007		;
assign memory[	567	]=	16'd	25040		;
assign memory[	568	]=	16'd	25072		;
assign memory[	569	]=	16'd	25105	     ;
assign memory[	570	]=	16'd	25137		;
assign memory[	571	]=	16'd	25169		;
assign memory[	572	]=	16'd	25201		;
assign memory[	573	]=	16'd	25233		;
assign memory[	574	]=	16'd	25265		;
assign memory[	575	]=	16'd	25297		;
assign memory[	576	]=	16'd	25329		;
assign memory[	577	]=	16'd	25361		;
assign memory[	578	]=	16'd	25393		;
assign memory[	579	]=	16'd	25425		;
assign memory[	580	]=	16'd	25456		;
assign memory[	581	]=	16'd	25488		;
assign memory[	582	]=	16'd	25519		;
assign memory[	583	]=	16'd	25551		;
assign memory[	584	]=	16'd	25582		;
assign memory[	585	]=	16'd	25614		;
assign memory[	586	]=	16'd	25645		;
assign memory[	587	]=	16'd	25676		;
assign memory[	588	]=	16'd	25708		;
assign memory[	589	]=	16'd	25739	     ;
assign memory[	590	]=	16'd	25770		;
assign memory[	591	]=	16'd	25801		;
assign memory[	592	]=	16'd	25832		;
assign memory[	593	]=	16'd	25863		;
assign memory[	594	]=	16'd	25893		;
assign memory[	595	]=	16'd	25924	     ;
assign memory[	596	]=	16'd	25955		;
assign memory[	597	]=	16'd	25986	     ;
assign memory[	598	]=	16'd	26016		;
assign memory[	599	]=	16'd	26047		;
assign memory[	600	]=	16'd	26077		;
assign memory[	601	]=	16'd	26108	     ;
assign memory[	602	]=	16'd	26138		;
assign memory[	603	]=	16'd	26168		;
assign memory[	604	]=	16'd	26198		;
assign memory[	605	]=	16'd	26229		;
assign memory[	606	]=	16'd	26259		;
assign memory[	607	]=	16'd	26289		;
assign memory[	608	]=	16'd	26319		;
assign memory[	609	]=	16'd	26349		;
assign memory[	610	]=	16'd	26378		;
assign memory[	611	]=	16'd	26408		;
assign memory[	612	]=	16'd	26438		;
assign memory[	613	]=	16'd	26468		;
assign memory[	614	]=	16'd	26497		;
assign memory[	615	]=	16'd	26527		;
assign memory[	616	]=	16'd	26556		;
assign memory[	617	]=	16'd	26586		;
assign memory[	618	]=	16'd	26615		;
assign memory[	619	]=	16'd	26644		;
assign memory[	620	]=	16'd	26674	     ;
assign memory[	621	]=	16'd	26703		;
assign memory[	622	]=	16'd	26732		;
assign memory[	623	]=	16'd	26761		;
assign memory[	624	]=	16'd	26790		;
assign memory[	625	]=	16'd	26819	     ;
assign memory[	626	]=	16'd	26848	     ;
assign memory[	627	]=	16'd	26876		;
assign memory[	628	]=	16'd	26905		;
assign memory[	629	]=	16'd	26934		;
assign memory[	630	]=	16'd	26962		;
assign memory[	631	]=	16'd	26991		;
assign memory[	632	]=	16'd	27019		;
assign memory[	633	]=	16'd	27048		;
assign memory[	634	]=	16'd	27076		;
assign memory[	635	]=	16'd	27104		;
assign memory[	636	]=	16'd	27133		;
assign memory[	637	]=	16'd	27161		;
assign memory[	638	]=	16'd	27189		;
assign memory[	639	]=	16'd	27217	     ;
assign memory[	640	]=	16'd	27245		;
assign memory[	641	]=	16'd	27273		;
assign memory[	642	]=	16'd	27300		;
assign memory[	643	]=	16'd	27328		;
assign memory[	644	]=	16'd	27356		;
assign memory[	645	]=	16'd	27384		;
assign memory[	646	]=	16'd	27411		;
assign memory[	647	]=	16'd	27439		;
assign memory[	648	]=	16'd	27466		;
assign memory[	649	]=	16'd	27493		;
assign memory[	650	]=	16'd	27521		;
assign memory[	651	]=	16'd	27548		;
assign memory[	652	]=	16'd	27575		;
assign memory[	653	]=	16'd	27602	     ;
assign memory[	654	]=	16'd	27629	     ;
assign memory[	655	]=	16'd	27656		;
assign memory[	656	]=	16'd	27683		;
assign memory[	657	]=	16'd	27710		;
assign memory[	658	]=	16'd	27737		;
assign memory[	659	]=	16'd	27764		;
assign memory[	660	]=	16'd	27790		;
assign memory[	661	]=	16'd	27817		;
assign memory[	662	]=	16'd	27843		;
assign memory[	663	]=	16'd	27870		;
assign memory[	664	]=	16'd	27896		;
assign memory[	665	]=	16'd	27923		;
assign memory[	666	]=	16'd	27949		;
assign memory[	667	]=	16'd	27975		;
assign memory[	668	]=	16'd	28001		;
assign memory[	669	]=	16'd	28027		;
assign memory[	670	]=	16'd	28053		;
assign memory[	671	]=	16'd	28079		;
assign memory[	672	]=	16'd	28105	     ;
assign memory[	673	]=	16'd	28131		;
assign memory[	674	]=	16'd	28157		;
assign memory[	675	]=	16'd	28182	     ;
assign memory[	676	]=	16'd	28208		;
assign memory[	677	]=	16'd	28234		;
assign memory[	678	]=	16'd	28259		;
assign memory[	679	]=	16'd	28284		;
assign memory[	680	]=	16'd	28310		;
assign memory[	681	]=	16'd	28335		;
assign memory[	682	]=	16'd	28360		;
assign memory[	683	]=	16'd	28385		;
assign memory[	684	]=	16'd	28411		;
assign memory[	685	]=	16'd	28436		;
assign memory[	686	]=	16'd	28460		;
assign memory[	687	]=	16'd	28485		;
assign memory[	688	]=	16'd	28510		;
assign memory[	689	]=	16'd	28535		;
assign memory[	690	]=	16'd	28560		;
assign memory[	691	]=	16'd	28584		;
assign memory[	692	]=	16'd	28609		;
assign memory[	693	]=	16'd	28633		;
assign memory[	694	]=	16'd	28658		;
assign memory[	695	]=	16'd	28682		;
assign memory[	696	]=	16'd	28706		;
assign memory[	697	]=	16'd	28730		;
assign memory[	698	]=	16'd	28755	     ;
assign memory[	699	]=	16'd	28779		;
assign memory[	700	]=	16'd	28803		;
assign memory[	701	]=	16'd	28827		;
assign memory[	702	]=	16'd	28850		;
assign memory[	703	]=	16'd	28874		;
assign memory[	704	]=	16'd	28898		;
assign memory[	705	]=	16'd	28922	     ;
assign memory[	706	]=	16'd	28945		;
assign memory[	707	]=	16'd	28969		;
assign memory[	708	]=	16'd	28992		;
assign memory[	709	]=	16'd	29016		;
assign memory[	710	]=	16'd	29039	     ;
assign memory[	711	]=	16'd	29062		;
assign memory[	712	]=	16'd	29085	     ;
assign memory[	713	]=	16'd	29108		;
assign memory[	714	]=	16'd	29131		;
assign memory[	715	]=	16'd	29154		;
assign memory[	716	]=	16'd	29177		;
assign memory[	717	]=	16'd	29200		;
assign memory[	718	]=	16'd	29223		;
assign memory[	719	]=	16'd	29246		;
assign memory[	720	]=	16'd	29268		;
assign memory[	721	]=	16'd	29291		;
assign memory[	722	]=	16'd	29313		;
assign memory[	723	]=	16'd	29336		;
assign memory[	724	]=	16'd	29358	     ;
assign memory[	725	]=	16'd	29380	     ;
assign memory[	726	]=	16'd	29403		;
assign memory[	727	]=	16'd	29425	     ;
assign memory[	728	]=	16'd	29447		;
assign memory[	729	]=	16'd	29469		;
assign memory[	730	]=	16'd	29491		;
assign memory[	731	]=	16'd	29513		;
assign memory[	732	]=	16'd	29534		;
assign memory[	733	]=	16'd	29556		;
assign memory[	734	]=	16'd	29578		;
assign memory[	735	]=	16'd	29599		;
assign memory[	736	]=	16'd	29621		;
assign memory[	737	]=	16'd	29642		;
assign memory[	738	]=	16'd	29664		;
assign memory[	739	]=	16'd	29685		;
assign memory[	740	]=	16'd	29706		;
assign memory[	741	]=	16'd	29728		;
assign memory[	742	]=	16'd	29749		;
assign memory[	743	]=	16'd	29770		;
assign memory[	744	]=	16'd	29791		;
assign memory[	745	]=	16'd	29812		;
assign memory[	746	]=	16'd	29832		;
assign memory[	747	]=	16'd	29853		;
assign memory[	748	]=	16'd	29874		;
assign memory[	749	]=	16'd	29894		;
assign memory[	750	]=	16'd	29915	     ;
assign memory[	751	]=	16'd	29936		;
assign memory[	752	]=	16'd	29956		;
assign memory[	753	]=	16'd	29976		;
assign memory[	754	]=	16'd	29997		;
assign memory[	755	]=	16'd	30017		;
assign memory[	756	]=	16'd	30037	     ;
assign memory[	757	]=	16'd	30057		;
assign memory[	758	]=	16'd	30077		;
assign memory[	759	]=	16'd	30097		;
assign memory[	760	]=	16'd	30117		;
assign memory[	761	]=	16'd	30136		;
assign memory[	762	]=	16'd	30156		;
assign memory[	763	]=	16'd	30176		;
assign memory[	764	]=	16'd	30195		;
assign memory[	765	]=	16'd	30215		;
assign memory[	766	]=	16'd	30234		;
assign memory[	767	]=	16'd	30253		;
assign memory[	768	]=	16'd	30273		;
assign memory[	769	]=	16'd	30292		;
assign memory[	770	]=	16'd	30311		;
assign memory[	771	]=	16'd	30330		;
assign memory[	772	]=	16'd	30349		;
assign memory[	773	]=	16'd	30368		;
assign memory[	774	]=	16'd	30387		;
assign memory[	775	]=	16'd	30406		;
assign memory[	776	]=	16'd	30424	     ;
assign memory[	777	]=	16'd	30443		;
assign memory[	778	]=	16'd	30462		;
assign memory[	779	]=	16'd	30480		;
assign memory[	780	]=	16'd	30498		;
assign memory[	781	]=	16'd	30517		;
assign memory[	782	]=	16'd	30535		;
assign memory[	783	]=	16'd	30553		;
assign memory[	784	]=	16'd	30571		;
assign memory[	785	]=	16'd	30589		;
assign memory[	786	]=	16'd	30607	     ;
assign memory[	787	]=	16'd	30625	     ;
assign memory[	788	]=	16'd	30643	     ;
assign memory[	789	]=	16'd	30661		;
assign memory[	790	]=	16'd	30679		;
assign memory[	791	]=	16'd	30696		;
assign memory[	792	]=	16'd	30714		;
assign memory[	793	]=	16'd	30731		;
assign memory[	794	]=	16'd	30749		;
assign memory[	795	]=	16'd	30766		;
assign memory[	796	]=	16'd	30783		;
assign memory[	797	]=	16'd	30800		;
assign memory[	798	]=	16'd	30818		;
assign memory[	799	]=	16'd	30835		;
assign memory[	800	]=	16'd	30852		;
assign memory[	801	]=	16'd	30868	     ;
assign memory[	802	]=	16'd	30885		;
assign memory[	803	]=	16'd	30902		;
assign memory[	804	]=	16'd	30919		;
assign memory[	805	]=	16'd	30935		;
assign memory[	806	]=	16'd	30952		;
assign memory[	807	]=	16'd	30968		;
assign memory[	808	]=	16'd	30985		;
assign memory[	809	]=	16'd	31001		;
assign memory[	810	]=	16'd	31017		;
assign memory[	811	]=	16'd	31033		;
assign memory[	812	]=	16'd	31050		;
assign memory[	813	]=	16'd	31066		;
assign memory[	814	]=	16'd	31082	     ;
assign memory[	815	]=	16'd	31097		;
assign memory[	816	]=	16'd	31113		;
assign memory[	817	]=	16'd	31129		;
assign memory[	818	]=	16'd	31145		;
assign memory[	819	]=	16'd	31160		;
assign memory[	820	]=	16'd	31176		;
assign memory[	821	]=	16'd	31191		;
assign memory[	822	]=	16'd	31206		;
assign memory[	823	]=	16'd	31222		;
assign memory[	824	]=	16'd	31237	     ;
assign memory[	825	]=	16'd	31252	     ;
assign memory[	826	]=	16'd	31267		;
assign memory[	827	]=	16'd	31282		;
assign memory[	828	]=	16'd	31297		;
assign memory[	829	]=	16'd	31312		;
assign memory[	830	]=	16'd	31327		;
assign memory[	831	]=	16'd	31341		;
assign memory[	832	]=	16'd	31356		;
assign memory[	833	]=	16'd	31371		;
assign memory[	834	]=	16'd	31385		;
assign memory[	835	]=	16'd	31400		;
assign memory[	836	]=	16'd	31414		;
assign memory[	837	]=	16'd	31428		;
assign memory[	838	]=	16'd	31442		;
assign memory[	839	]=	16'd	31456		;
assign memory[	840	]=	16'd	31470		;
assign memory[	841	]=	16'd	31484		;
assign memory[	842	]=	16'd	31498		;
assign memory[	843	]=	16'd	31512		;
assign memory[	844	]=	16'd	31526		;
assign memory[	845	]=	16'd	31539		;
assign memory[	846	]=	16'd	31553		;
assign memory[	847	]=	16'd	31567	     ;
assign memory[	848	]=	16'd	31580		;
assign memory[	849	]=	16'd	31593		;
assign memory[	850	]=	16'd	31607		;
assign memory[	851	]=	16'd	31620		;
assign memory[	852	]=	16'd	31633		;
assign memory[	853	]=	16'd	31646		;
assign memory[	854	]=	16'd	31659		;
assign memory[	855	]=	16'd	31672		;
assign memory[	856	]=	16'd	31685		;
assign memory[	857	]=	16'd	31698		;
assign memory[	858	]=	16'd	31710		;
assign memory[	859	]=	16'd	31723		;
assign memory[	860	]=	16'd	31736		;
assign memory[	861	]=	16'd	31748		;
assign memory[	862	]=	16'd	31760		;
assign memory[	863	]=	16'd	31773		;
assign memory[	864	]=	16'd	31785		;
assign memory[	865	]=	16'd	31797		;
assign memory[	866	]=	16'd	31809		;
assign memory[	867	]=	16'd	31821		;
assign memory[	868	]=	16'd	31833		;
assign memory[	869	]=	16'd	31845		;
assign memory[	870	]=	16'd	31857		;
assign memory[	871	]=	16'd	31869		;
assign memory[	872	]=	16'd	31880		;
assign memory[	873	]=	16'd	31892		;
assign memory[	874	]=	16'd	31903	     ;
assign memory[	875	]=	16'd	31915		;
assign memory[	876	]=	16'd	31926		;
assign memory[	877	]=	16'd	31937		;
assign memory[	878	]=	16'd	31949		;
assign memory[	879	]=	16'd	31960		;
assign memory[	880	]=	16'd	31971	     ;
assign memory[	881	]=	16'd	31982		;
assign memory[	882	]=	16'd	31993		;
assign memory[	883	]=	16'd	32004		;
assign memory[	884	]=	16'd	32014		;
assign memory[	885	]=	16'd	32025	     ;
assign memory[	886	]=	16'd	32036		;
assign memory[	887	]=	16'd	32046		;
assign memory[	888	]=	16'd	32057		;
assign memory[	889	]=	16'd	32067		;
assign memory[	890	]=	16'd	32077		;
assign memory[	891	]=	16'd	32087		;
assign memory[	892	]=	16'd	32098		;
assign memory[	893	]=	16'd	32108		;
assign memory[	894	]=	16'd	32118		;
assign memory[	895	]=	16'd	32128		;
assign memory[	896	]=	16'd	32137	     ;
assign memory[	897	]=	16'd	32147		;
assign memory[	898	]=	16'd	32157		;
assign memory[	899	]=	16'd	32166		;
assign memory[	900	]=	16'd	32176		;
assign memory[	901	]=	16'd	32185		;
assign memory[	902	]=	16'd	32195		;
assign memory[	903	]=	16'd	32204		;
assign memory[	904	]=	16'd	32213		;
assign memory[	905	]=	16'd	32223	     ;
assign memory[	906	]=	16'd	32232		;
assign memory[	907	]=	16'd	32241		;
assign memory[	908	]=	16'd	32250		;
assign memory[	909	]=	16'd	32258		;
assign memory[	910	]=	16'd	32267		;
assign memory[	911	]=	16'd	32276		;
assign memory[	912	]=	16'd	32285		;
assign memory[	913	]=	16'd	32293		;
assign memory[	914	]=	16'd	32302		;
assign memory[	915	]=	16'd	32310		;
assign memory[	916	]=	16'd	32318		;
assign memory[	917	]=	16'd	32327	     ;
assign memory[	918	]=	16'd	32335		;
assign memory[	919	]=	16'd	32343		;
assign memory[	920	]=	16'd	32351		;
assign memory[	921	]=	16'd	32359		;
assign memory[	922	]=	16'd	32367		;
assign memory[	923	]=	16'd	32375		;
assign memory[	924	]=	16'd	32382		;
assign memory[	925	]=	16'd	32390		;
assign memory[	926	]=	16'd	32397		;
assign memory[	927	]=	16'd	32405		;
assign memory[	928	]=	16'd	32412	     ;
assign memory[	929	]=	16'd	32420		;
assign memory[	930	]=	16'd	32427		;
assign memory[	931	]=	16'd	32434		;
assign memory[	932	]=	16'd	32441	     ;
assign memory[	933	]=	16'd	32448		;
assign memory[	934	]=	16'd	32455		;
assign memory[	935	]=	16'd	32462		;
assign memory[	936	]=	16'd	32469		;
assign memory[	937	]=	16'd	32476		;
assign memory[	938	]=	16'd	32482	     ;
assign memory[	939	]=	16'd	32489		;
assign memory[	940	]=	16'd	32495		;
assign memory[	941	]=	16'd	32502	     ;
assign memory[	942	]=	16'd	32508		;
assign memory[	943	]=	16'd	32514		;
assign memory[	944	]=	16'd	32521		;
assign memory[	945	]=	16'd	32527		;
assign memory[	946	]=	16'd	32533		;
assign memory[	947	]=	16'd	32539	     ;
assign memory[	948	]=	16'd	32545		;
assign memory[	949	]=	16'd	32550		;
assign memory[	950	]=	16'd	32556		;
assign memory[	951	]=	16'd	32562		;
assign memory[	952	]=	16'd	32567	     ;
assign memory[	953	]=	16'd	32573		;
assign memory[	954	]=	16'd	32578		;
assign memory[	955	]=	16'd	32584	     ;
assign memory[	956	]=	16'd	32589		;
assign memory[	957	]=	16'd	32594		;
assign memory[	958	]=	16'd	32599		;
assign memory[	959	]=	16'd	32604		;
assign memory[	960	]=	16'd	32609		;
assign memory[	961	]=	16'd	32614		;
assign memory[	962	]=	16'd	32619		;
assign memory[	963	]=	16'd	32624		;
assign memory[	964	]=	16'd	32628		;
assign memory[	965	]=	16'd	32633		;
assign memory[	966	]=	16'd	32637		;
assign memory[	967	]=	16'd	32642		;
assign memory[	968	]=	16'd	32646		;
assign memory[	969	]=	16'd	32650		;
assign memory[	970	]=	16'd	32655		;
assign memory[	971	]=	16'd	32659		;
assign memory[	972	]=	16'd	32663		;
assign memory[	973	]=	16'd	32667		;
assign memory[	974	]=	16'd	32671	     ;
assign memory[	975	]=	16'd	32674		;
assign memory[	976	]=	16'd	32678		;
assign memory[	977	]=	16'd	32682	     ;
assign memory[	978	]=	16'd	32685		;
assign memory[	979	]=	16'd	32689		;
assign memory[	980	]=	16'd	32692		;
assign memory[	981	]=	16'd	32696	     ;
assign memory[	982	]=	16'd	32699		;
assign memory[	983	]=	16'd	32702		;
assign memory[	984	]=	16'd	32705		;
assign memory[	985	]=	16'd	32708		;
assign memory[	986	]=	16'd	32711		;
assign memory[	987	]=	16'd	32714		;
assign memory[	988	]=	16'd	32717		;
assign memory[	989	]=	16'd	32720		;
assign memory[	990	]=	16'd	32722		;
assign memory[	991	]=	16'd	32725		;
assign memory[	992	]=	16'd	32728		;
assign memory[	993	]=	16'd	32730	     ;
assign memory[	994	]=	16'd	32732		;
assign memory[	995	]=	16'd	32735		;
assign memory[	996	]=	16'd	32737		;
assign memory[	997	]=	16'd	32739		;
assign memory[	998	]=	16'd	32741		;
assign memory[	999	]=	16'd	32743		;
assign memory[	1000	]=	16'd	32745		;
assign memory[	1001	]=	16'd	32747	     ;
assign memory[	1002	]=	16'd	32748		;
assign memory[	1003	]=	16'd	32750		;
assign memory[	1004	]=	16'd	32752		;
assign memory[	1005	]=	16'd	32753		;
assign memory[	1006	]=	16'd	32755		;
assign memory[	1007	]=	16'd	32756		;
assign memory[	1008	]=	16'd	32757		;
assign memory[	1009	]=	16'd	32758		;
assign memory[	1010	]=	16'd	32759		;
assign memory[	1011	]=	16'd	32760	     ;
assign memory[	1012	]=	16'd	32761		;
assign memory[	1013	]=	16'd	32762		;
assign memory[	1014	]=	16'd	32763		;
assign memory[	1015	]=	16'd	32764		;
assign memory[	1016	]=	16'd	32765		;
assign memory[	1017	]=	16'd	32765	     ;
assign memory[	1018	]=	16'd	32766		;
assign memory[	1019	]=	16'd	32766		;
assign memory[	1020	]=	16'd	32766		;
assign memory[	1021	]=	16'd	32767		;
assign memory[	1022	]=	16'd	32767		;
assign memory[	1023	]=	16'd	32767		;

endmodule
