library verilog;
use verilog.vl_types.all;
entity song_reader_tb_v is
    generic(
        delay           : integer := 10
    );
end song_reader_tb_v;
