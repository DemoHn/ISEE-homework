library verilog;
use verilog.vl_types.all;
entity music_player_tb_v is
    generic(
        delay           : integer := 10
    );
end music_player_tb_v;
